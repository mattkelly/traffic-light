TODO placeholder for testbench for overall system
