TODO placeholder for overall system with TMR
